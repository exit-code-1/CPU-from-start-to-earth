`define IF_TO_ID_WD 33
`define ID_TO_EX_WD 163
`define EX_TO_MEM_WD 82
`define MEM_TO_WB_WD 70
`define BR_WD 33
`define DATA_SRAM_WD 69
`define WB_TO_RF_WD 38
`define EX_TO_ID_WD 44
`define MEM_TO_ID_WD 38
`define ID_TO_PC_WD 33
`define INIT 32'h00000000
`define StallBus 6
`define NoStop 1'b0
`define Stop 1'b1
`define DELAY_TO_EX_WD 33
`define SW 6'b101011
`define SB 6'b101000
`define SH 6'b101001
`define SWL 6'b101010
`define SWR 6'b101100
`define LB 6'b101011
`define LBU 6'b101011
`define LW 6'b100011
